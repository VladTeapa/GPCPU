localparam logic [7:0] ROM_STICK_0[255:0] = '{
0:8'h3b, 1:8'h00, 2:8'h42, 3:8'h00, 4:8'h00, 5:8'h30, 6:8'h41, 7:8'h40, 8:8'h02, 9:8'h48, 
10:8'h10, 11:8'h58, 12:8'h10, 13:8'h42, 14:8'h00, 15:8'h00, 16:8'h01, 17:8'h16, 18:8'h10, 19:8'h74, 
20:8'h00, 21:8'h17, 22:8'h70, 23:8'h00, 24:8'h00, 25:8'h16, 26:8'h17, 27:8'h14, 28:8'h41, 29:8'h00, 
30:8'h0a, 31:8'h10, 32:8'h13, 33:8'h12, 34:8'h41, 35:8'hc0, 36:8'h02, 37:8'h41, 38:8'h40, 39:8'h06, 
40:8'h43, 41:8'h50, 42:8'h41, 43:8'h40, 44:8'h09, 45:8'h43, 46:8'h60, 47:8'h1c, 48:8'hfe, 49:8'h75, 
50:8'h05, 51:8'h00, 52:8'h01, 53:8'h02, 54:8'h03, 55:8'h04, 56:8'h05, 57:8'h06, 58:8'h07, 59:8'h08, 
60:8'h09, default:8'h00
};
